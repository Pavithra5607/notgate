module not_gate_dataflow (input a,
                          output y);
  assign y = ~a;
endmodule